/*
	Port_ID Decoder
	
	Project: III Digitales
	Designer: Luis Leon
	Developer: Luis Leon
	Start Date: 13-Oct-2016
	End Date: -- No yet --
	Description: This is the port id decoder for selecting the output of the controller
*/

module Port_ID_Decoder(
		input [7:0] Port_ID,
		output reg[1:0] DataSelect
	);
	
	always @*
	begin
		begin
			case(Port_ID)
			8'h01: DataSelect = 2'd0;
			8'h02: DataSelect = 2'd1;
			8'h03: DataSelect = 2'd2;
			default: DataSelect = 2'd3;
			endcase
		end
	
	end

endmodule