`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    17:37:47 10/16/2016 
// Design Name: 
// Module Name:    deco_id 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module deco_id(id_port, actRTC, actVGA, actTeclado, actsonido, dir);
	input[7:0] id_port;
	output actRTC, actVGA, actTeclado, actsonido;
	output [7:0] dir;
	reg actRTC, actVGA, actTeclado, actsonido;
	reg [7:0] dir;
	always @ *
	begin
		case (id_port)
		8'd1:
		begin
			actRTC=1;
			actVGA=0; 
			actTeclado=0; 
			actsonido=0;
			dir=8'd0;
		end
		8'd2:
		begin
			actRTC=1;
			actVGA=0; 
			actTeclado=0; 
			actsonido=0;
			dir=8'd1;
		end
		8'd3:
		begin
			actRTC=1;
			actVGA=0; 
			actTeclado=0; 
			actsonido=0;
			dir=8'd2;
		end
		8'd4:
		begin
			actRTC=1;
			actVGA=0; 
			actTeclado=0; 
			actsonido=0;
			dir=8'hF0;
		end
		8'd5:
		begin
			actRTC=0;
			actVGA=0; 
			actTeclado=1; 
			actsonido=0;
			dir=8'd1;
		end
		8'd6:
		begin
			actRTC=0;
			actVGA=0; 
			actTeclado=1; 
			actsonido=0;
			dir=8'd2;
		end
		8'd7:
		begin
			actRTC=0;
			actVGA=0; 
			actTeclado=1; 
			actsonido=0;
			dir=8'd3;
		end
		8'd11:
		begin
			actRTC=1;
			actVGA=0; 
			actTeclado=0; 
			actsonido=0;
			dir=8'd11;
		end
		//segundos
		8'd17:
		begin
			actRTC=1;
			actVGA=0; 
			actTeclado=0; 
			actsonido=0;
			dir=8'd33;
		end
		//minutos
		8'd18:
		begin
			actRTC=1;
			actVGA=0; 
			actTeclado=0; 
			actsonido=0;
			dir=8'd34;
		end
		//horas
		8'd19:
		begin
			actRTC=1;
			actVGA=0; 
			actTeclado=0; 
			actsonido=0;
			dir=8'd35;
		end
		//dias
		8'd20:
		begin
			actRTC=1;
			actVGA=0; 
			actTeclado=0; 
			actsonido=0;
			dir=8'd36;
		end
		//meses
		8'd21:
		begin
			actRTC=1;
			actVGA=0; 
			actTeclado=0; 
			actsonido=0;
			dir=8'd37;
		end
		//year
		8'd22:
		begin
			actRTC=1;
			actVGA=0; 
			actTeclado=0; 
			actsonido=0;
			dir=8'd38;
		end
		//segundos timer
		8'd23:
		begin
			actRTC=1;
			actVGA=0; 
			actTeclado=0; 
			actsonido=0;
			dir=8'h41;
		end
		//minutos timer
		8'd24:
		begin
			actRTC=1;
			actVGA=0; 
			actTeclado=0; 
			actsonido=0;
			dir=8'h42;
		end
		//horas timer
		8'd25:
		begin
			actRTC=1;
			actVGA=0; 
			actTeclado=0; 
			actsonido=0;
			dir=8'h43;
		end
		8'd26:
		begin
			actRTC=1;
			actVGA=0; 
			actTeclado=0; 
			actsonido=0;
			dir=8'd10;
		end
		//puntero
		8'd27:
		begin
			actRTC=1;
			actVGA=0; 
			actTeclado=0; 
			actsonido=0;
			dir=8'd11;
		end
		//timer activado
		8'd28:
		begin
			actRTC=1;
			actVGA=0; 
			actTeclado=0; 
			actsonido=0;
			dir=8'd12;
		end
		8'd40:
		begin
			actRTC=0;
			actVGA=1; 
			actTeclado=0; 
			actsonido=0;
			dir=8'd40;
		end
		8'd41:
		begin
			actRTC=0;
			actVGA=1; 
			actTeclado=0; 
			actsonido=0;
			dir=8'd41;
		end
		8'd42:
		begin
			actRTC=0;
			actVGA=1; 
			actTeclado=0; 
			actsonido=0;
			dir=8'd42;
		end
		8'd43:
		begin
			actRTC=0;
			actVGA=1; 
			actTeclado=0; 
			actsonido=0;
			dir=8'd45;
		end
		8'd44:
		begin
			actRTC=0;
			actVGA=1; 
			actTeclado=0; 
			actsonido=0;
			dir=8'd44;
		end
		8'd45:
		begin
			actRTC=0;
			actVGA=1; 
			actTeclado=0; 
			actsonido=0;
			dir=8'd43;
		end
		8'd46:
		begin
			actRTC=0;
			actVGA=1; 
			actTeclado=0; 
			actsonido=0;
			dir=8'd46;
		end
		8'd47:
		begin
			actRTC=0;
			actVGA=1; 
			actTeclado=0; 
			actsonido=0;
			dir=8'd47;
		end
		8'd48:
		begin
			actRTC=0;
			actVGA=1; 
			actTeclado=0; 
			actsonido=0;
			dir=8'd48;
		end
		8'd49:
		begin
			actRTC=0;
			actVGA=1; 
			actTeclado=0; 
			actsonido=0;
			dir=8'd49;
		end
		8'd51:
		begin
			actRTC=0;
			actVGA=1; 
			actTeclado=0; 
			actsonido=0;
			dir=8'd51;
		end
		8'd50:
		begin
			actRTC=0;
			actVGA=1; 
			actTeclado=0; 
			actsonido=0;
			dir=8'd50;
		end
		default:
		begin
			actRTC=0;
			actVGA=0; 
			actTeclado=0; 
			actsonido=0;
			dir=8'd0;
		end
		endcase
	end
endmodule
